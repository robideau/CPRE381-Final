 -- adder.vhd
 --
 -- The adders used for calculating PC-plus-4 and branch targets
 -- CprE 381
 --
 -- Zhao Zhang, Fall 2013
 --

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.mips32.all;

entity adder is
  generic (DELAY : time := 19.0 ns);
  port (src1    : in  m32_word;
        src2    : in  m32_word;
        result  : out m32_word);
end entity;

-- Behavior modeling of ADDER
architecture behavior of adder is
begin
  ADD : process (src1, src2)
    variable a : integer;
    variable b : integer;
    variable c : integer;
  begin
    -- Pre-calculate
    a := to_integer(signed(src1));
    b := to_integer(signed(src2));
    c := a + b;
    
    -- Convert integer to 32-bit signal
    result <= std_logic_vector(to_signed(c, result'length)) after DELAY;
  end process;
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.mips32.all;

entity adder_structural is
   port (src1    : in  m32_word;
        src2    : in  m32_word;
        result  : out m32_word);
end entity;

architecture structural of adder_structural is

component full_adder
  port (i_x0  : in std_logic;
       i_x1  : in std_logic;
       i_C  : in std_logic;
       o_Co : out std_logic;
       o_Y  : out std_logic); 
end component;

signal c_out : std_logic_vector(31 downto 0);

begin

Adder_0 : full_adder
port map(
    i_x0 => src1(0),
    i_x1 => src2(0),
    i_C => '0',
    o_Co => c_out(0),
    o_Y => result(0)
  );

G1: for i in 1 to 31 generate
  Adder_i : full_adder
    port map(
      i_x0 => src1(i),
      i_x1 => src2(i),
      i_C => c_out(i-1),
      o_Co => c_out(i),
      o_Y => result(i)
    );
  end generate;
end structural;